module MUX4_1(inA, inB, inC, inD, sel);
input 
